module bola(

);

endmodule