module cursor(
    input clk,
    input [5:0] size,
    input draw,
    input [10:0] x,
    input [10:0] y,
    input z

  // complemente seus sinais aqui
);

endmodule

