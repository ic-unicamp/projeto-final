module tela(
    input CLOCK_50,
    input reset,
    input [9:0] BordaBarraX,
    input [9:0] BordaBarraY,
    input [9:0] LarguraBarra, 
    input [9:0] AlturaBarra, 
    input [9:0] BolaNaveX,  
    input [9:0] BolaNaveY,
    input [9:0] BolaInimigaX,
    input [9:0] BolaInimigaY,
    input [9:0] LadoBola,
    output reg [7:0] VGA_R,    
    output reg [7:0] VGA_G, 
    output reg [7:0] VGA_B, 
    output wire VGA_HS,  
    output wire VGA_VS,
    output wire VGA_BLANK_N,
    output wire VGA_SYNC_N, 
	output wire VGA_CLK, 
	input perdeu
);  
    wire [9:0] VGA_X;
    wire [9:0] VGA_Y; 
    wire ativo;
    reg [0:3071] texto = 3072'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111011111010001011111000011111010001011111011111000000000000001000001000101101101000000001000101000101000001000100000000000000101110111110101010111110000100010100010111110111110000000000000010001010001010001010000000010001001010010000010010000000000000001111101000101000101111100001111100010001111101000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	 reg xTela = 0;
	 reg yTela = 0;
	 reg [4:0] inicio;
	 reg [32:0] indice;
	 
	vga v(
		.CLOCK_50(CLOCK_50),
		.reset(reset),
		.VGA_CLK(VGA_CLK),
        .VGA_HS(VGA_HS),
        .VGA_VS(VGA_VS),
        .VGA_BLANK_N(VGA_BLANK_N),
        .VGA_SYNC_N(VGA_SYNC_N),
		.x(VGA_X),
		.y(VGA_Y),
		.ativo(ativo)
	);

    always @(posedge CLOCK_50 or posedge reset) begin // implementar a lógica que será usada para "imprimir" na tela
        if (reset) begin
		   	VGA_R = 0;
            VGA_G = 0;
            VGA_B = 0;
        end else begin
            if (ativo && !perdeu) begin
                if ((BordaBarraX + 144 <= VGA_X ) && (VGA_X <= 144 + BordaBarraX + LarguraBarra) && 
                    (BordaBarraY + 35 <= VGA_Y) && (VGA_Y <= BordaBarraY + 35 + AlturaBarra)) begin // da barra
                    VGA_R = 255;
                    VGA_G = 255;
                    VGA_B = 255;
                    end else if ((BolaX + 144 <= VGA_X ) && (VGA_X <= 144 + BolaX + LadoBola) && 
                        (BolaY + 35 <= VGA_Y) && (VGA_Y <= BolaY + 35 + LadoBola)) begin //o da bola
                    VGA_R = 255;
                    VGA_G = 255;
                    VGA_B = 255;
                end else begin
                    VGA_R = 0; 
                    VGA_G = 50;
                    VGA_B = 50;
                end
				end else if (ativo && perdeu) begin
                    indice = (VGA_Y - 35) / 10 * (64) + ((VGA_X - 144) / 10); 
                    if (texto[indice] == 1) begin
                        VGA_R = 255;
                        VGA_G = 255;
                        VGA_B = 255;
                    end else begin
                        VGA_R = 255;
                        VGA_G = 0;
                        VGA_B = 0;                   
                    end
				
            end else begin 
                    VGA_R = 0;
                    VGA_G = 0;
                    VGA_B = 0;  
                    indice = 0;
            end
        end
    end

endmodule