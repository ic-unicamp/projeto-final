module projeto(

);

endmodule